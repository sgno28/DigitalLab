`include "pc.sv"
`include "rom.sv"

module instruction_memory (
    input CLK, reset
)